--  C:\USERS\DICKOVER\DOCUMENTS\...\EVBD_MAIN_FIFO.vhd
--  VHDL code created by Xilinx's StateCAD 10.1
--  Mon Mar 21 18:16:17 2016

--  This VHDL code (for use with Xilinx XST) was generated using: 
--  enumerated state assignment with structured code format.
--  Minimization is enabled,  implied else is enabled, 
--  and outputs are area optimized.

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY EVBD_MAIN_FIFO IS
	PORT (CLK,A_GO,A_Trailer,B_GO,B_Trailer,Block_Done,EVEN,Event_Done,
		Event_Trig_Go,RESET_N: IN std_logic;
		A_SEL,aevbd_rd_en,B_SEL,bevbd_rd_en,Block_Header_Go1,Block_Header_Go2,
			Block_Trail_GO1,Block_Trail_GO2,Clear_chip_ev,DEC_Evt_Trig_cnt,
			Filler_Word_GO1,Filler_Word_GO2,FWEN_N,INC_chip_ev,INC_Event_cnt,word_cnt : 
			OUT std_logic);
END;

ARCHITECTURE BEHAVIOR OF EVBD_MAIN_FIFO IS
	TYPE type_sreg IS (Block_Done_S,Block_Header1,Block_Header2,Block_Trailer1,
		Block_Trailer2,Choose_A,Choose_B,ehold,End_Event,Event_Done_S,Filler_Word1,
		Filler_Word2,idle,Inc_A,INC_B,Start,STATE0,STATE1,STATE2,STATE3,STATE4,STATE5
		,STATE6,STATE7,STATE8,STATE9,STATE10,STATE11,STATE12,STATE13,STATE14,STATE15,
		STATE16);
	SIGNAL sreg, next_sreg : type_sreg;
BEGIN
	PROCESS (CLK, next_sreg)
	BEGIN
		IF CLK='1' AND CLK'event THEN
			sreg <= next_sreg;
		END IF;
	END PROCESS;

	PROCESS (sreg,A_GO,A_Trailer,B_GO,B_Trailer,Block_Done,EVEN,Event_Done,
		Event_Trig_Go,RESET_N)
	BEGIN
		A_SEL <= '0'; aevbd_rd_en <= '0'; B_SEL <= '0'; bevbd_rd_en <= '0'; 
			Block_Header_Go1 <= '0'; Block_Header_Go2 <= '0'; Block_Trail_GO1 <= '0'; 
			Block_Trail_GO2 <= '0'; Clear_chip_ev <= '0'; DEC_Evt_Trig_cnt <= '0'; 
			Filler_Word_GO1 <= '0'; Filler_Word_GO2 <= '0'; FWEN_N <= '0'; INC_chip_ev <=
			 '0'; INC_Event_cnt <= '0'; word_cnt <= '0'; 

		next_sreg<=Block_Done_S;

		IF ( RESET_N='0' ) THEN
			next_sreg<=idle;
			A_SEL<='0';
			aevbd_rd_en<='0';
			B_SEL<='0';
			bevbd_rd_en<='0';
			Block_Header_Go1<='0';
			Block_Header_Go2<='0';
			Block_Trail_GO1<='0';
			Block_Trail_GO2<='0';
			Clear_chip_ev<='0';
			DEC_Evt_Trig_cnt<='0';
			Filler_Word_GO1<='0';
			Filler_Word_GO2<='0';
			FWEN_N<='0';
			INC_chip_ev<='0';
			INC_Event_cnt<='0';
			word_cnt<='0';
		ELSE
			CASE sreg IS
				WHEN Block_Done_S =>
					A_SEL<='0';
					aevbd_rd_en<='0';
					B_SEL<='0';
					bevbd_rd_en<='0';
					Block_Header_Go1<='0';
					Block_Header_Go2<='0';
					Block_Trail_GO1<='0';
					Block_Trail_GO2<='0';
					Clear_chip_ev<='0';
					DEC_Evt_Trig_cnt<='0';
					Filler_Word_GO1<='0';
					Filler_Word_GO2<='0';
					FWEN_N<='0';
					INC_chip_ev<='0';
					INC_Event_cnt<='0';
					word_cnt<='0';
					IF ( EVEN='1' ) THEN
						next_sreg<=Filler_Word1;
					END IF;
					IF ( EVEN='0' ) THEN
						next_sreg<=Block_Trailer1;
					END IF;
				WHEN Block_Header1 =>
					A_SEL<='0';
					aevbd_rd_en<='0';
					B_SEL<='0';
					bevbd_rd_en<='0';
					Block_Header_Go2<='0';
					Block_Trail_GO1<='0';
					Block_Trail_GO2<='0';
					Clear_chip_ev<='0';
					DEC_Evt_Trig_cnt<='0';
					Filler_Word_GO1<='0';
					Filler_Word_GO2<='0';
					INC_chip_ev<='0';
					INC_Event_cnt<='0';
					Block_Header_Go1<='1';
					FWEN_N<='1';
					word_cnt<='1';
					next_sreg<=Block_Header2;
				WHEN Block_Header2 =>
					A_SEL<='0';
					aevbd_rd_en<='0';
					B_SEL<='0';
					bevbd_rd_en<='0';
					Block_Header_Go1<='0';
					Block_Trail_GO1<='0';
					Block_Trail_GO2<='0';
					Clear_chip_ev<='0';
					DEC_Evt_Trig_cnt<='0';
					Filler_Word_GO1<='0';
					Filler_Word_GO2<='0';
					INC_chip_ev<='0';
					INC_Event_cnt<='0';
					Block_Header_Go2<='1';
					FWEN_N<='1';
					word_cnt<='1';
					next_sreg<=Start;
				WHEN Block_Trailer1 =>
					A_SEL<='0';
					aevbd_rd_en<='0';
					B_SEL<='0';
					bevbd_rd_en<='0';
					Block_Header_Go1<='0';
					Block_Header_Go2<='0';
					Block_Trail_GO2<='0';
					Clear_chip_ev<='0';
					DEC_Evt_Trig_cnt<='0';
					Filler_Word_GO1<='0';
					Filler_Word_GO2<='0';
					INC_chip_ev<='0';
					INC_Event_cnt<='0';
					Block_Trail_GO1<='1';
					FWEN_N<='1';
					word_cnt<='1';
					next_sreg<=Block_Trailer2;
				WHEN Block_Trailer2 =>
					A_SEL<='0';
					aevbd_rd_en<='0';
					B_SEL<='0';
					bevbd_rd_en<='0';
					Block_Header_Go1<='0';
					Block_Header_Go2<='0';
					Block_Trail_GO1<='0';
					Clear_chip_ev<='0';
					DEC_Evt_Trig_cnt<='0';
					Filler_Word_GO1<='0';
					Filler_Word_GO2<='0';
					INC_chip_ev<='0';
					INC_Event_cnt<='0';
					Block_Trail_GO2<='1';
					FWEN_N<='1';
					word_cnt<='1';
					next_sreg<=STATE3;
				WHEN Choose_A =>
					B_SEL<='0';
					bevbd_rd_en<='0';
					Block_Header_Go1<='0';
					Block_Header_Go2<='0';
					Block_Trail_GO1<='0';
					Block_Trail_GO2<='0';
					Clear_chip_ev<='0';
					DEC_Evt_Trig_cnt<='0';
					Filler_Word_GO1<='0';
					Filler_Word_GO2<='0';
					INC_chip_ev<='0';
					INC_Event_cnt<='0';
					A_SEL<='1';
					aevbd_rd_en<='1';
					FWEN_N<='1';
					word_cnt<='1';
					IF ( A_Trailer='1' ) THEN
						next_sreg<=Inc_A;
					 ELSE
						next_sreg<=Choose_A;
					END IF;
				WHEN Choose_B =>
					A_SEL<='0';
					aevbd_rd_en<='0';
					Block_Header_Go1<='0';
					Block_Header_Go2<='0';
					Block_Trail_GO1<='0';
					Block_Trail_GO2<='0';
					Clear_chip_ev<='0';
					DEC_Evt_Trig_cnt<='0';
					Filler_Word_GO1<='0';
					Filler_Word_GO2<='0';
					INC_chip_ev<='0';
					INC_Event_cnt<='0';
					B_SEL<='1';
					bevbd_rd_en<='1';
					FWEN_N<='1';
					word_cnt<='1';
					IF ( B_Trailer='1' ) THEN
						next_sreg<=INC_B;
					 ELSE
						next_sreg<=Choose_B;
					END IF;
				WHEN ehold =>
					A_SEL<='0';
					aevbd_rd_en<='0';
					B_SEL<='0';
					bevbd_rd_en<='0';
					Block_Header_Go1<='0';
					Block_Header_Go2<='0';
					Block_Trail_GO1<='0';
					Block_Trail_GO2<='0';
					Clear_chip_ev<='0';
					DEC_Evt_Trig_cnt<='0';
					Filler_Word_GO1<='0';
					Filler_Word_GO2<='0';
					FWEN_N<='0';
					INC_chip_ev<='0';
					INC_Event_cnt<='0';
					word_cnt<='0';
					next_sreg<=End_Event;
				WHEN End_Event =>
					A_SEL<='0';
					aevbd_rd_en<='0';
					B_SEL<='0';
					bevbd_rd_en<='0';
					Block_Header_Go1<='0';
					Block_Header_Go2<='0';
					Block_Trail_GO1<='0';
					Block_Trail_GO2<='0';
					Clear_chip_ev<='0';
					DEC_Evt_Trig_cnt<='0';
					Filler_Word_GO1<='0';
					Filler_Word_GO2<='0';
					FWEN_N<='0';
					INC_chip_ev<='0';
					INC_Event_cnt<='0';
					word_cnt<='0';
					IF ( Block_Done='1' ) THEN
						next_sreg<=Block_Done_S;
					ELSIF ( Block_Done='0' ) THEN
						next_sreg<=Start;
					END IF;
				WHEN Event_Done_S =>
					A_SEL<='0';
					aevbd_rd_en<='0';
					B_SEL<='0';
					bevbd_rd_en<='0';
					Block_Header_Go1<='0';
					Block_Header_Go2<='0';
					Block_Trail_GO1<='0';
					Block_Trail_GO2<='0';
					Filler_Word_GO1<='0';
					Filler_Word_GO2<='0';
					FWEN_N<='0';
					INC_chip_ev<='0';
					word_cnt<='0';
					INC_Event_cnt<='1';
					DEC_Evt_Trig_cnt<='1';
					Clear_chip_ev<='1';
					next_sreg<=ehold;
				WHEN Filler_Word1 =>
					A_SEL<='0';
					aevbd_rd_en<='0';
					B_SEL<='0';
					bevbd_rd_en<='0';
					Block_Header_Go1<='0';
					Block_Header_Go2<='0';
					Block_Trail_GO1<='0';
					Block_Trail_GO2<='0';
					Clear_chip_ev<='0';
					DEC_Evt_Trig_cnt<='0';
					Filler_Word_GO2<='0';
					INC_chip_ev<='0';
					INC_Event_cnt<='0';
					Filler_Word_GO1<='1';
					FWEN_N<='1';
					word_cnt<='1';
					next_sreg<=Filler_Word2;
				WHEN Filler_Word2 =>
					A_SEL<='0';
					aevbd_rd_en<='0';
					B_SEL<='0';
					bevbd_rd_en<='0';
					Block_Header_Go1<='0';
					Block_Header_Go2<='0';
					Block_Trail_GO1<='0';
					Block_Trail_GO2<='0';
					Clear_chip_ev<='0';
					DEC_Evt_Trig_cnt<='0';
					Filler_Word_GO1<='0';
					INC_chip_ev<='0';
					INC_Event_cnt<='0';
					Filler_Word_GO2<='1';
					FWEN_N<='1';
					word_cnt<='1';
					next_sreg<=Block_Trailer1;
				WHEN idle =>
					A_SEL<='0';
					aevbd_rd_en<='0';
					B_SEL<='0';
					bevbd_rd_en<='0';
					Block_Header_Go1<='0';
					Block_Header_Go2<='0';
					Block_Trail_GO1<='0';
					Block_Trail_GO2<='0';
					Clear_chip_ev<='0';
					DEC_Evt_Trig_cnt<='0';
					Filler_Word_GO1<='0';
					Filler_Word_GO2<='0';
					FWEN_N<='0';
					INC_chip_ev<='0';
					INC_Event_cnt<='0';
					word_cnt<='0';
					next_sreg<=STATE7;
				WHEN Inc_A =>
					aevbd_rd_en<='0';
					B_SEL<='0';
					bevbd_rd_en<='0';
					Block_Header_Go1<='0';
					Block_Header_Go2<='0';
					Block_Trail_GO1<='0';
					Block_Trail_GO2<='0';
					Clear_chip_ev<='0';
					DEC_Evt_Trig_cnt<='0';
					Filler_Word_GO1<='0';
					Filler_Word_GO2<='0';
					INC_Event_cnt<='0';
					A_SEL<='1';
					FWEN_N<='1';
					word_cnt<='1';
					INC_chip_ev<='1';
					next_sreg<=STATE2;
				WHEN INC_B =>
					A_SEL<='0';
					aevbd_rd_en<='0';
					bevbd_rd_en<='0';
					Block_Header_Go1<='0';
					Block_Header_Go2<='0';
					Block_Trail_GO1<='0';
					Block_Trail_GO2<='0';
					Clear_chip_ev<='0';
					DEC_Evt_Trig_cnt<='0';
					Filler_Word_GO1<='0';
					Filler_Word_GO2<='0';
					INC_Event_cnt<='0';
					B_SEL<='1';
					FWEN_N<='1';
					word_cnt<='1';
					INC_chip_ev<='1';
					next_sreg<=STATE1;
				WHEN Start =>
					A_SEL<='0';
					aevbd_rd_en<='0';
					B_SEL<='0';
					bevbd_rd_en<='0';
					Block_Header_Go1<='0';
					Block_Header_Go2<='0';
					Block_Trail_GO1<='0';
					Block_Trail_GO2<='0';
					Clear_chip_ev<='0';
					DEC_Evt_Trig_cnt<='0';
					Filler_Word_GO1<='0';
					Filler_Word_GO2<='0';
					FWEN_N<='0';
					INC_chip_ev<='0';
					INC_Event_cnt<='0';
					word_cnt<='0';
					IF ( A_GO='1' ) THEN
						next_sreg<=STATE13;
					ELSIF ( B_GO='1' ) THEN
						next_sreg<=STATE15;
					ELSIF ( Event_Done='1' ) THEN
						next_sreg<=Event_Done_S;
					 ELSE
						next_sreg<=Start;
					END IF;
				WHEN STATE0 =>
					A_SEL<='0';
					aevbd_rd_en<='0';
					B_SEL<='0';
					bevbd_rd_en<='0';
					Block_Header_Go1<='0';
					Block_Header_Go2<='0';
					Block_Trail_GO1<='0';
					Block_Trail_GO2<='0';
					Clear_chip_ev<='0';
					DEC_Evt_Trig_cnt<='0';
					Filler_Word_GO1<='0';
					Filler_Word_GO2<='0';
					FWEN_N<='0';
					INC_chip_ev<='0';
					INC_Event_cnt<='0';
					word_cnt<='0';
					next_sreg<=idle;
				WHEN STATE1 =>
					A_SEL<='0';
					aevbd_rd_en<='0';
					bevbd_rd_en<='0';
					Block_Header_Go1<='0';
					Block_Header_Go2<='0';
					Block_Trail_GO1<='0';
					Block_Trail_GO2<='0';
					Clear_chip_ev<='0';
					DEC_Evt_Trig_cnt<='0';
					Filler_Word_GO1<='0';
					Filler_Word_GO2<='0';
					FWEN_N<='0';
					INC_chip_ev<='0';
					INC_Event_cnt<='0';
					word_cnt<='0';
					B_SEL<='1';
					next_sreg<=Start;
				WHEN STATE2 =>
					aevbd_rd_en<='0';
					B_SEL<='0';
					bevbd_rd_en<='0';
					Block_Header_Go1<='0';
					Block_Header_Go2<='0';
					Block_Trail_GO1<='0';
					Block_Trail_GO2<='0';
					Clear_chip_ev<='0';
					DEC_Evt_Trig_cnt<='0';
					Filler_Word_GO1<='0';
					Filler_Word_GO2<='0';
					FWEN_N<='0';
					INC_chip_ev<='0';
					INC_Event_cnt<='0';
					word_cnt<='0';
					A_SEL<='1';
					next_sreg<=Start;
				WHEN STATE3 =>
					A_SEL<='0';
					aevbd_rd_en<='0';
					B_SEL<='0';
					bevbd_rd_en<='0';
					Block_Header_Go1<='0';
					Block_Header_Go2<='0';
					Block_Trail_GO1<='0';
					Block_Trail_GO2<='0';
					Clear_chip_ev<='0';
					DEC_Evt_Trig_cnt<='0';
					Filler_Word_GO1<='0';
					Filler_Word_GO2<='0';
					FWEN_N<='0';
					INC_chip_ev<='0';
					INC_Event_cnt<='0';
					word_cnt<='0';
					next_sreg<=STATE4;
				WHEN STATE4 =>
					A_SEL<='0';
					aevbd_rd_en<='0';
					B_SEL<='0';
					bevbd_rd_en<='0';
					Block_Header_Go1<='0';
					Block_Header_Go2<='0';
					Block_Trail_GO1<='0';
					Block_Trail_GO2<='0';
					Clear_chip_ev<='0';
					DEC_Evt_Trig_cnt<='0';
					Filler_Word_GO1<='0';
					Filler_Word_GO2<='0';
					FWEN_N<='0';
					INC_chip_ev<='0';
					INC_Event_cnt<='0';
					word_cnt<='0';
					next_sreg<=STATE8;
				WHEN STATE5 =>
					B_SEL<='0';
					bevbd_rd_en<='0';
					Block_Header_Go1<='0';
					Block_Header_Go2<='0';
					Block_Trail_GO1<='0';
					Block_Trail_GO2<='0';
					Clear_chip_ev<='0';
					DEC_Evt_Trig_cnt<='0';
					Filler_Word_GO1<='0';
					Filler_Word_GO2<='0';
					FWEN_N<='0';
					INC_chip_ev<='0';
					INC_Event_cnt<='0';
					word_cnt<='0';
					A_SEL<='1';
					aevbd_rd_en<='1';
					next_sreg<=Choose_A;
				WHEN STATE6 =>
					A_SEL<='0';
					aevbd_rd_en<='0';
					Block_Header_Go1<='0';
					Block_Header_Go2<='0';
					Block_Trail_GO1<='0';
					Block_Trail_GO2<='0';
					Clear_chip_ev<='0';
					DEC_Evt_Trig_cnt<='0';
					Filler_Word_GO1<='0';
					Filler_Word_GO2<='0';
					FWEN_N<='0';
					INC_chip_ev<='0';
					INC_Event_cnt<='0';
					word_cnt<='0';
					B_SEL<='1';
					bevbd_rd_en<='1';
					next_sreg<=Choose_B;
				WHEN STATE7 =>
					A_SEL<='0';
					aevbd_rd_en<='0';
					B_SEL<='0';
					bevbd_rd_en<='0';
					Block_Header_Go1<='0';
					Block_Header_Go2<='0';
					Block_Trail_GO1<='0';
					Block_Trail_GO2<='0';
					Clear_chip_ev<='0';
					DEC_Evt_Trig_cnt<='0';
					Filler_Word_GO1<='0';
					Filler_Word_GO2<='0';
					FWEN_N<='0';
					INC_chip_ev<='0';
					INC_Event_cnt<='0';
					word_cnt<='0';
					next_sreg<=STATE12;
				WHEN STATE8 =>
					A_SEL<='0';
					aevbd_rd_en<='0';
					B_SEL<='0';
					bevbd_rd_en<='0';
					Block_Header_Go1<='0';
					Block_Header_Go2<='0';
					Block_Trail_GO1<='0';
					Block_Trail_GO2<='0';
					Clear_chip_ev<='0';
					DEC_Evt_Trig_cnt<='0';
					Filler_Word_GO1<='0';
					Filler_Word_GO2<='0';
					FWEN_N<='0';
					INC_chip_ev<='0';
					INC_Event_cnt<='0';
					word_cnt<='0';
					next_sreg<=STATE0;
				WHEN STATE9 =>
					A_SEL<='0';
					aevbd_rd_en<='0';
					B_SEL<='0';
					bevbd_rd_en<='0';
					Block_Header_Go1<='0';
					Block_Header_Go2<='0';
					Block_Trail_GO1<='0';
					Block_Trail_GO2<='0';
					Clear_chip_ev<='0';
					DEC_Evt_Trig_cnt<='0';
					Filler_Word_GO1<='0';
					Filler_Word_GO2<='0';
					FWEN_N<='0';
					INC_chip_ev<='0';
					INC_Event_cnt<='0';
					word_cnt<='0';
					next_sreg<=STATE10;
				WHEN STATE10 =>
					A_SEL<='0';
					aevbd_rd_en<='0';
					B_SEL<='0';
					bevbd_rd_en<='0';
					Block_Header_Go1<='0';
					Block_Header_Go2<='0';
					Block_Trail_GO1<='0';
					Block_Trail_GO2<='0';
					Clear_chip_ev<='0';
					DEC_Evt_Trig_cnt<='0';
					Filler_Word_GO1<='0';
					Filler_Word_GO2<='0';
					FWEN_N<='0';
					INC_chip_ev<='0';
					INC_Event_cnt<='0';
					word_cnt<='0';
					next_sreg<=STATE11;
				WHEN STATE11 =>
					A_SEL<='0';
					aevbd_rd_en<='0';
					B_SEL<='0';
					bevbd_rd_en<='0';
					Block_Header_Go1<='0';
					Block_Header_Go2<='0';
					Block_Trail_GO1<='0';
					Block_Trail_GO2<='0';
					Clear_chip_ev<='0';
					DEC_Evt_Trig_cnt<='0';
					Filler_Word_GO1<='0';
					Filler_Word_GO2<='0';
					FWEN_N<='0';
					INC_chip_ev<='0';
					INC_Event_cnt<='0';
					word_cnt<='0';
					IF ( Event_Trig_Go='1' ) THEN
						next_sreg<=Block_Header1;
					 ELSE
						next_sreg<=STATE11;
					END IF;
				WHEN STATE12 =>
					A_SEL<='0';
					aevbd_rd_en<='0';
					B_SEL<='0';
					bevbd_rd_en<='0';
					Block_Header_Go1<='0';
					Block_Header_Go2<='0';
					Block_Trail_GO1<='0';
					Block_Trail_GO2<='0';
					Clear_chip_ev<='0';
					DEC_Evt_Trig_cnt<='0';
					Filler_Word_GO1<='0';
					Filler_Word_GO2<='0';
					FWEN_N<='0';
					INC_chip_ev<='0';
					INC_Event_cnt<='0';
					word_cnt<='0';
					next_sreg<=STATE9;
				WHEN STATE13 =>
					A_SEL<='0';
					aevbd_rd_en<='0';
					B_SEL<='0';
					bevbd_rd_en<='0';
					Block_Header_Go1<='0';
					Block_Header_Go2<='0';
					Block_Trail_GO1<='0';
					Block_Trail_GO2<='0';
					Clear_chip_ev<='0';
					DEC_Evt_Trig_cnt<='0';
					Filler_Word_GO1<='0';
					Filler_Word_GO2<='0';
					FWEN_N<='0';
					INC_chip_ev<='0';
					INC_Event_cnt<='0';
					word_cnt<='0';
					next_sreg<=STATE14;
				WHEN STATE14 =>
					A_SEL<='0';
					aevbd_rd_en<='0';
					B_SEL<='0';
					bevbd_rd_en<='0';
					Block_Header_Go1<='0';
					Block_Header_Go2<='0';
					Block_Trail_GO1<='0';
					Block_Trail_GO2<='0';
					Clear_chip_ev<='0';
					DEC_Evt_Trig_cnt<='0';
					Filler_Word_GO1<='0';
					Filler_Word_GO2<='0';
					FWEN_N<='0';
					INC_chip_ev<='0';
					INC_Event_cnt<='0';
					word_cnt<='0';
					next_sreg<=STATE5;
				WHEN STATE15 =>
					A_SEL<='0';
					aevbd_rd_en<='0';
					B_SEL<='0';
					bevbd_rd_en<='0';
					Block_Header_Go1<='0';
					Block_Header_Go2<='0';
					Block_Trail_GO1<='0';
					Block_Trail_GO2<='0';
					Clear_chip_ev<='0';
					DEC_Evt_Trig_cnt<='0';
					Filler_Word_GO1<='0';
					Filler_Word_GO2<='0';
					FWEN_N<='0';
					INC_chip_ev<='0';
					INC_Event_cnt<='0';
					word_cnt<='0';
					next_sreg<=STATE16;
				WHEN STATE16 =>
					A_SEL<='0';
					aevbd_rd_en<='0';
					B_SEL<='0';
					bevbd_rd_en<='0';
					Block_Header_Go1<='0';
					Block_Header_Go2<='0';
					Block_Trail_GO1<='0';
					Block_Trail_GO2<='0';
					Clear_chip_ev<='0';
					DEC_Evt_Trig_cnt<='0';
					Filler_Word_GO1<='0';
					Filler_Word_GO2<='0';
					FWEN_N<='0';
					INC_chip_ev<='0';
					INC_Event_cnt<='0';
					word_cnt<='0';
					next_sreg<=STATE6;
				WHEN OTHERS =>
			END CASE;
		END IF;
	END PROCESS;
END BEHAVIOR;
